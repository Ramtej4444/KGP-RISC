`timescale 1ns / 1ps

module ADD( input [31:0] in_0,
				input [31:0] in_1,
				output [31:0] out
    );
	
assign out = in_0 + in_1;


endmodule
